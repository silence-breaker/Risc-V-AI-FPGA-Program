package my_types_pkg;
  typedef enum logic [1:0] {
    W_ZERO = 2'b00,
    W_POS  = 2'b01,
    W_NEG  = 2'b11
  } tern_t;
endpackage
